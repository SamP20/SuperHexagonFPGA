library verilog;
use verilog.vl_types.all;
entity random_gen_tb is
end random_gen_tb;
