// Lookup table for generating sin and cos values
module sincos(
	input clk,
	input [9:0]angle,
	output reg signed [11:0]sin,
	output reg signed [11:0]cos
);

reg signed [11:0]lookup[0:1023];

always @(posedge clk) begin
	sin <= lookup[angle];
	cos <= lookup[angle+10'd256];
end

initial begin
	lookup[0] = 12'sd0;
	lookup[1] = 12'sd12;
	lookup[2] = 12'sd25;
	lookup[3] = 12'sd37;
	lookup[4] = 12'sd50;
	lookup[5] = 12'sd62;
	lookup[6] = 12'sd75;
	lookup[7] = 12'sd87;
	lookup[8] = 12'sd100;
	lookup[9] = 12'sd113;
	lookup[10] = 12'sd125;
	lookup[11] = 12'sd138;
	lookup[12] = 12'sd150;
	lookup[13] = 12'sd163;
	lookup[14] = 12'sd175;
	lookup[15] = 12'sd188;
	lookup[16] = 12'sd200;
	lookup[17] = 12'sd213;
	lookup[18] = 12'sd225;
	lookup[19] = 12'sd238;
	lookup[20] = 12'sd250;
	lookup[21] = 12'sd263;
	lookup[22] = 12'sd275;
	lookup[23] = 12'sd288;
	lookup[24] = 12'sd300;
	lookup[25] = 12'sd312;
	lookup[26] = 12'sd325;
	lookup[27] = 12'sd337;
	lookup[28] = 12'sd350;
	lookup[29] = 12'sd362;
	lookup[30] = 12'sd374;
	lookup[31] = 12'sd387;
	lookup[32] = 12'sd399;
	lookup[33] = 12'sd411;
	lookup[34] = 12'sd424;
	lookup[35] = 12'sd436;
	lookup[36] = 12'sd448;
	lookup[37] = 12'sd460;
	lookup[38] = 12'sd473;
	lookup[39] = 12'sd485;
	lookup[40] = 12'sd497;
	lookup[41] = 12'sd509;
	lookup[42] = 12'sd521;
	lookup[43] = 12'sd534;
	lookup[44] = 12'sd546;
	lookup[45] = 12'sd558;
	lookup[46] = 12'sd570;
	lookup[47] = 12'sd582;
	lookup[48] = 12'sd594;
	lookup[49] = 12'sd606;
	lookup[50] = 12'sd618;
	lookup[51] = 12'sd630;
	lookup[52] = 12'sd642;
	lookup[53] = 12'sd654;
	lookup[54] = 12'sd666;
	lookup[55] = 12'sd678;
	lookup[56] = 12'sd689;
	lookup[57] = 12'sd701;
	lookup[58] = 12'sd713;
	lookup[59] = 12'sd725;
	lookup[60] = 12'sd737;
	lookup[61] = 12'sd748;
	lookup[62] = 12'sd760;
	lookup[63] = 12'sd772;
	lookup[64] = 12'sd783;
	lookup[65] = 12'sd795;
	lookup[66] = 12'sd806;
	lookup[67] = 12'sd818;
	lookup[68] = 12'sd829;
	lookup[69] = 12'sd841;
	lookup[70] = 12'sd852;
	lookup[71] = 12'sd864;
	lookup[72] = 12'sd875;
	lookup[73] = 12'sd886;
	lookup[74] = 12'sd898;
	lookup[75] = 12'sd909;
	lookup[76] = 12'sd920;
	lookup[77] = 12'sd932;
	lookup[78] = 12'sd943;
	lookup[79] = 12'sd954;
	lookup[80] = 12'sd965;
	lookup[81] = 12'sd976;
	lookup[82] = 12'sd987;
	lookup[83] = 12'sd998;
	lookup[84] = 12'sd1009;
	lookup[85] = 12'sd1020;
	lookup[86] = 12'sd1031;
	lookup[87] = 12'sd1042;
	lookup[88] = 12'sd1052;
	lookup[89] = 12'sd1063;
	lookup[90] = 12'sd1074;
	lookup[91] = 12'sd1085;
	lookup[92] = 12'sd1095;
	lookup[93] = 12'sd1106;
	lookup[94] = 12'sd1116;
	lookup[95] = 12'sd1127;
	lookup[96] = 12'sd1137;
	lookup[97] = 12'sd1148;
	lookup[98] = 12'sd1158;
	lookup[99] = 12'sd1168;
	lookup[100] = 12'sd1179;
	lookup[101] = 12'sd1189;
	lookup[102] = 12'sd1199;
	lookup[103] = 12'sd1209;
	lookup[104] = 12'sd1219;
	lookup[105] = 12'sd1230;
	lookup[106] = 12'sd1240;
	lookup[107] = 12'sd1250;
	lookup[108] = 12'sd1259;
	lookup[109] = 12'sd1269;
	lookup[110] = 12'sd1279;
	lookup[111] = 12'sd1289;
	lookup[112] = 12'sd1299;
	lookup[113] = 12'sd1308;
	lookup[114] = 12'sd1318;
	lookup[115] = 12'sd1328;
	lookup[116] = 12'sd1337;
	lookup[117] = 12'sd1347;
	lookup[118] = 12'sd1356;
	lookup[119] = 12'sd1366;
	lookup[120] = 12'sd1375;
	lookup[121] = 12'sd1384;
	lookup[122] = 12'sd1393;
	lookup[123] = 12'sd1403;
	lookup[124] = 12'sd1412;
	lookup[125] = 12'sd1421;
	lookup[126] = 12'sd1430;
	lookup[127] = 12'sd1439;
	lookup[128] = 12'sd1448;
	lookup[129] = 12'sd1457;
	lookup[130] = 12'sd1465;
	lookup[131] = 12'sd1474;
	lookup[132] = 12'sd1483;
	lookup[133] = 12'sd1491;
	lookup[134] = 12'sd1500;
	lookup[135] = 12'sd1509;
	lookup[136] = 12'sd1517;
	lookup[137] = 12'sd1525;
	lookup[138] = 12'sd1534;
	lookup[139] = 12'sd1542;
	lookup[140] = 12'sd1550;
	lookup[141] = 12'sd1558;
	lookup[142] = 12'sd1567;
	lookup[143] = 12'sd1575;
	lookup[144] = 12'sd1583;
	lookup[145] = 12'sd1591;
	lookup[146] = 12'sd1598;
	lookup[147] = 12'sd1606;
	lookup[148] = 12'sd1614;
	lookup[149] = 12'sd1622;
	lookup[150] = 12'sd1629;
	lookup[151] = 12'sd1637;
	lookup[152] = 12'sd1644;
	lookup[153] = 12'sd1652;
	lookup[154] = 12'sd1659;
	lookup[155] = 12'sd1667;
	lookup[156] = 12'sd1674;
	lookup[157] = 12'sd1681;
	lookup[158] = 12'sd1688;
	lookup[159] = 12'sd1695;
	lookup[160] = 12'sd1702;
	lookup[161] = 12'sd1709;
	lookup[162] = 12'sd1716;
	lookup[163] = 12'sd1723;
	lookup[164] = 12'sd1730;
	lookup[165] = 12'sd1736;
	lookup[166] = 12'sd1743;
	lookup[167] = 12'sd1750;
	lookup[168] = 12'sd1756;
	lookup[169] = 12'sd1763;
	lookup[170] = 12'sd1769;
	lookup[171] = 12'sd1775;
	lookup[172] = 12'sd1781;
	lookup[173] = 12'sd1788;
	lookup[174] = 12'sd1794;
	lookup[175] = 12'sd1800;
	lookup[176] = 12'sd1806;
	lookup[177] = 12'sd1812;
	lookup[178] = 12'sd1817;
	lookup[179] = 12'sd1823;
	lookup[180] = 12'sd1829;
	lookup[181] = 12'sd1834;
	lookup[182] = 12'sd1840;
	lookup[183] = 12'sd1845;
	lookup[184] = 12'sd1851;
	lookup[185] = 12'sd1856;
	lookup[186] = 12'sd1861;
	lookup[187] = 12'sd1867;
	lookup[188] = 12'sd1872;
	lookup[189] = 12'sd1877;
	lookup[190] = 12'sd1882;
	lookup[191] = 12'sd1887;
	lookup[192] = 12'sd1892;
	lookup[193] = 12'sd1896;
	lookup[194] = 12'sd1901;
	lookup[195] = 12'sd1906;
	lookup[196] = 12'sd1910;
	lookup[197] = 12'sd1915;
	lookup[198] = 12'sd1919;
	lookup[199] = 12'sd1924;
	lookup[200] = 12'sd1928;
	lookup[201] = 12'sd1932;
	lookup[202] = 12'sd1936;
	lookup[203] = 12'sd1940;
	lookup[204] = 12'sd1944;
	lookup[205] = 12'sd1948;
	lookup[206] = 12'sd1952;
	lookup[207] = 12'sd1956;
	lookup[208] = 12'sd1959;
	lookup[209] = 12'sd1963;
	lookup[210] = 12'sd1966;
	lookup[211] = 12'sd1970;
	lookup[212] = 12'sd1973;
	lookup[213] = 12'sd1977;
	lookup[214] = 12'sd1980;
	lookup[215] = 12'sd1983;
	lookup[216] = 12'sd1986;
	lookup[217] = 12'sd1989;
	lookup[218] = 12'sd1992;
	lookup[219] = 12'sd1995;
	lookup[220] = 12'sd1998;
	lookup[221] = 12'sd2000;
	lookup[222] = 12'sd2003;
	lookup[223] = 12'sd2006;
	lookup[224] = 12'sd2008;
	lookup[225] = 12'sd2011;
	lookup[226] = 12'sd2013;
	lookup[227] = 12'sd2015;
	lookup[228] = 12'sd2017;
	lookup[229] = 12'sd2019;
	lookup[230] = 12'sd2021;
	lookup[231] = 12'sd2023;
	lookup[232] = 12'sd2025;
	lookup[233] = 12'sd2027;
	lookup[234] = 12'sd2029;
	lookup[235] = 12'sd2031;
	lookup[236] = 12'sd2032;
	lookup[237] = 12'sd2034;
	lookup[238] = 12'sd2035;
	lookup[239] = 12'sd2036;
	lookup[240] = 12'sd2038;
	lookup[241] = 12'sd2039;
	lookup[242] = 12'sd2040;
	lookup[243] = 12'sd2041;
	lookup[244] = 12'sd2042;
	lookup[245] = 12'sd2043;
	lookup[246] = 12'sd2044;
	lookup[247] = 12'sd2044;
	lookup[248] = 12'sd2045;
	lookup[249] = 12'sd2046;
	lookup[250] = 12'sd2046;
	lookup[251] = 12'sd2047;
	lookup[252] = 12'sd2047;
	lookup[253] = 12'sd2047;
	lookup[254] = 12'sd2047;
	lookup[255] = 12'sd2047;
	lookup[256] = 12'sd2047;
	lookup[257] = 12'sd2047;
	lookup[258] = 12'sd2047;
	lookup[259] = 12'sd2047;
	lookup[260] = 12'sd2047;
	lookup[261] = 12'sd2047;
	lookup[262] = 12'sd2046;
	lookup[263] = 12'sd2046;
	lookup[264] = 12'sd2045;
	lookup[265] = 12'sd2044;
	lookup[266] = 12'sd2044;
	lookup[267] = 12'sd2043;
	lookup[268] = 12'sd2042;
	lookup[269] = 12'sd2041;
	lookup[270] = 12'sd2040;
	lookup[271] = 12'sd2039;
	lookup[272] = 12'sd2038;
	lookup[273] = 12'sd2036;
	lookup[274] = 12'sd2035;
	lookup[275] = 12'sd2034;
	lookup[276] = 12'sd2032;
	lookup[277] = 12'sd2031;
	lookup[278] = 12'sd2029;
	lookup[279] = 12'sd2027;
	lookup[280] = 12'sd2025;
	lookup[281] = 12'sd2023;
	lookup[282] = 12'sd2021;
	lookup[283] = 12'sd2019;
	lookup[284] = 12'sd2017;
	lookup[285] = 12'sd2015;
	lookup[286] = 12'sd2013;
	lookup[287] = 12'sd2011;
	lookup[288] = 12'sd2008;
	lookup[289] = 12'sd2006;
	lookup[290] = 12'sd2003;
	lookup[291] = 12'sd2000;
	lookup[292] = 12'sd1998;
	lookup[293] = 12'sd1995;
	lookup[294] = 12'sd1992;
	lookup[295] = 12'sd1989;
	lookup[296] = 12'sd1986;
	lookup[297] = 12'sd1983;
	lookup[298] = 12'sd1980;
	lookup[299] = 12'sd1977;
	lookup[300] = 12'sd1973;
	lookup[301] = 12'sd1970;
	lookup[302] = 12'sd1966;
	lookup[303] = 12'sd1963;
	lookup[304] = 12'sd1959;
	lookup[305] = 12'sd1956;
	lookup[306] = 12'sd1952;
	lookup[307] = 12'sd1948;
	lookup[308] = 12'sd1944;
	lookup[309] = 12'sd1940;
	lookup[310] = 12'sd1936;
	lookup[311] = 12'sd1932;
	lookup[312] = 12'sd1928;
	lookup[313] = 12'sd1924;
	lookup[314] = 12'sd1919;
	lookup[315] = 12'sd1915;
	lookup[316] = 12'sd1910;
	lookup[317] = 12'sd1906;
	lookup[318] = 12'sd1901;
	lookup[319] = 12'sd1896;
	lookup[320] = 12'sd1892;
	lookup[321] = 12'sd1887;
	lookup[322] = 12'sd1882;
	lookup[323] = 12'sd1877;
	lookup[324] = 12'sd1872;
	lookup[325] = 12'sd1867;
	lookup[326] = 12'sd1861;
	lookup[327] = 12'sd1856;
	lookup[328] = 12'sd1851;
	lookup[329] = 12'sd1845;
	lookup[330] = 12'sd1840;
	lookup[331] = 12'sd1834;
	lookup[332] = 12'sd1829;
	lookup[333] = 12'sd1823;
	lookup[334] = 12'sd1817;
	lookup[335] = 12'sd1812;
	lookup[336] = 12'sd1806;
	lookup[337] = 12'sd1800;
	lookup[338] = 12'sd1794;
	lookup[339] = 12'sd1788;
	lookup[340] = 12'sd1781;
	lookup[341] = 12'sd1775;
	lookup[342] = 12'sd1769;
	lookup[343] = 12'sd1763;
	lookup[344] = 12'sd1756;
	lookup[345] = 12'sd1750;
	lookup[346] = 12'sd1743;
	lookup[347] = 12'sd1736;
	lookup[348] = 12'sd1730;
	lookup[349] = 12'sd1723;
	lookup[350] = 12'sd1716;
	lookup[351] = 12'sd1709;
	lookup[352] = 12'sd1702;
	lookup[353] = 12'sd1695;
	lookup[354] = 12'sd1688;
	lookup[355] = 12'sd1681;
	lookup[356] = 12'sd1674;
	lookup[357] = 12'sd1667;
	lookup[358] = 12'sd1659;
	lookup[359] = 12'sd1652;
	lookup[360] = 12'sd1644;
	lookup[361] = 12'sd1637;
	lookup[362] = 12'sd1629;
	lookup[363] = 12'sd1622;
	lookup[364] = 12'sd1614;
	lookup[365] = 12'sd1606;
	lookup[366] = 12'sd1598;
	lookup[367] = 12'sd1591;
	lookup[368] = 12'sd1583;
	lookup[369] = 12'sd1575;
	lookup[370] = 12'sd1567;
	lookup[371] = 12'sd1558;
	lookup[372] = 12'sd1550;
	lookup[373] = 12'sd1542;
	lookup[374] = 12'sd1534;
	lookup[375] = 12'sd1525;
	lookup[376] = 12'sd1517;
	lookup[377] = 12'sd1509;
	lookup[378] = 12'sd1500;
	lookup[379] = 12'sd1491;
	lookup[380] = 12'sd1483;
	lookup[381] = 12'sd1474;
	lookup[382] = 12'sd1465;
	lookup[383] = 12'sd1457;
	lookup[384] = 12'sd1448;
	lookup[385] = 12'sd1439;
	lookup[386] = 12'sd1430;
	lookup[387] = 12'sd1421;
	lookup[388] = 12'sd1412;
	lookup[389] = 12'sd1403;
	lookup[390] = 12'sd1393;
	lookup[391] = 12'sd1384;
	lookup[392] = 12'sd1375;
	lookup[393] = 12'sd1366;
	lookup[394] = 12'sd1356;
	lookup[395] = 12'sd1347;
	lookup[396] = 12'sd1337;
	lookup[397] = 12'sd1328;
	lookup[398] = 12'sd1318;
	lookup[399] = 12'sd1308;
	lookup[400] = 12'sd1299;
	lookup[401] = 12'sd1289;
	lookup[402] = 12'sd1279;
	lookup[403] = 12'sd1269;
	lookup[404] = 12'sd1259;
	lookup[405] = 12'sd1250;
	lookup[406] = 12'sd1240;
	lookup[407] = 12'sd1230;
	lookup[408] = 12'sd1219;
	lookup[409] = 12'sd1209;
	lookup[410] = 12'sd1199;
	lookup[411] = 12'sd1189;
	lookup[412] = 12'sd1179;
	lookup[413] = 12'sd1168;
	lookup[414] = 12'sd1158;
	lookup[415] = 12'sd1148;
	lookup[416] = 12'sd1137;
	lookup[417] = 12'sd1127;
	lookup[418] = 12'sd1116;
	lookup[419] = 12'sd1106;
	lookup[420] = 12'sd1095;
	lookup[421] = 12'sd1085;
	lookup[422] = 12'sd1074;
	lookup[423] = 12'sd1063;
	lookup[424] = 12'sd1052;
	lookup[425] = 12'sd1042;
	lookup[426] = 12'sd1031;
	lookup[427] = 12'sd1020;
	lookup[428] = 12'sd1009;
	lookup[429] = 12'sd998;
	lookup[430] = 12'sd987;
	lookup[431] = 12'sd976;
	lookup[432] = 12'sd965;
	lookup[433] = 12'sd954;
	lookup[434] = 12'sd943;
	lookup[435] = 12'sd932;
	lookup[436] = 12'sd920;
	lookup[437] = 12'sd909;
	lookup[438] = 12'sd898;
	lookup[439] = 12'sd886;
	lookup[440] = 12'sd875;
	lookup[441] = 12'sd864;
	lookup[442] = 12'sd852;
	lookup[443] = 12'sd841;
	lookup[444] = 12'sd829;
	lookup[445] = 12'sd818;
	lookup[446] = 12'sd806;
	lookup[447] = 12'sd795;
	lookup[448] = 12'sd783;
	lookup[449] = 12'sd772;
	lookup[450] = 12'sd760;
	lookup[451] = 12'sd748;
	lookup[452] = 12'sd737;
	lookup[453] = 12'sd725;
	lookup[454] = 12'sd713;
	lookup[455] = 12'sd701;
	lookup[456] = 12'sd689;
	lookup[457] = 12'sd678;
	lookup[458] = 12'sd666;
	lookup[459] = 12'sd654;
	lookup[460] = 12'sd642;
	lookup[461] = 12'sd630;
	lookup[462] = 12'sd618;
	lookup[463] = 12'sd606;
	lookup[464] = 12'sd594;
	lookup[465] = 12'sd582;
	lookup[466] = 12'sd570;
	lookup[467] = 12'sd558;
	lookup[468] = 12'sd546;
	lookup[469] = 12'sd534;
	lookup[470] = 12'sd521;
	lookup[471] = 12'sd509;
	lookup[472] = 12'sd497;
	lookup[473] = 12'sd485;
	lookup[474] = 12'sd473;
	lookup[475] = 12'sd460;
	lookup[476] = 12'sd448;
	lookup[477] = 12'sd436;
	lookup[478] = 12'sd424;
	lookup[479] = 12'sd411;
	lookup[480] = 12'sd399;
	lookup[481] = 12'sd387;
	lookup[482] = 12'sd374;
	lookup[483] = 12'sd362;
	lookup[484] = 12'sd350;
	lookup[485] = 12'sd337;
	lookup[486] = 12'sd325;
	lookup[487] = 12'sd312;
	lookup[488] = 12'sd300;
	lookup[489] = 12'sd288;
	lookup[490] = 12'sd275;
	lookup[491] = 12'sd263;
	lookup[492] = 12'sd250;
	lookup[493] = 12'sd238;
	lookup[494] = 12'sd225;
	lookup[495] = 12'sd213;
	lookup[496] = 12'sd200;
	lookup[497] = 12'sd188;
	lookup[498] = 12'sd175;
	lookup[499] = 12'sd163;
	lookup[500] = 12'sd150;
	lookup[501] = 12'sd138;
	lookup[502] = 12'sd125;
	lookup[503] = 12'sd113;
	lookup[504] = 12'sd100;
	lookup[505] = 12'sd87;
	lookup[506] = 12'sd75;
	lookup[507] = 12'sd62;
	lookup[508] = 12'sd50;
	lookup[509] = 12'sd37;
	lookup[510] = 12'sd25;
	lookup[511] = 12'sd12;
	lookup[512] = 12'sd0;
	lookup[513] = -12'sd12;
	lookup[514] = -12'sd25;
	lookup[515] = -12'sd37;
	lookup[516] = -12'sd50;
	lookup[517] = -12'sd62;
	lookup[518] = -12'sd75;
	lookup[519] = -12'sd87;
	lookup[520] = -12'sd100;
	lookup[521] = -12'sd113;
	lookup[522] = -12'sd125;
	lookup[523] = -12'sd138;
	lookup[524] = -12'sd150;
	lookup[525] = -12'sd163;
	lookup[526] = -12'sd175;
	lookup[527] = -12'sd188;
	lookup[528] = -12'sd200;
	lookup[529] = -12'sd213;
	lookup[530] = -12'sd225;
	lookup[531] = -12'sd238;
	lookup[532] = -12'sd250;
	lookup[533] = -12'sd263;
	lookup[534] = -12'sd275;
	lookup[535] = -12'sd288;
	lookup[536] = -12'sd300;
	lookup[537] = -12'sd312;
	lookup[538] = -12'sd325;
	lookup[539] = -12'sd337;
	lookup[540] = -12'sd350;
	lookup[541] = -12'sd362;
	lookup[542] = -12'sd374;
	lookup[543] = -12'sd387;
	lookup[544] = -12'sd399;
	lookup[545] = -12'sd411;
	lookup[546] = -12'sd424;
	lookup[547] = -12'sd436;
	lookup[548] = -12'sd448;
	lookup[549] = -12'sd460;
	lookup[550] = -12'sd473;
	lookup[551] = -12'sd485;
	lookup[552] = -12'sd497;
	lookup[553] = -12'sd509;
	lookup[554] = -12'sd521;
	lookup[555] = -12'sd534;
	lookup[556] = -12'sd546;
	lookup[557] = -12'sd558;
	lookup[558] = -12'sd570;
	lookup[559] = -12'sd582;
	lookup[560] = -12'sd594;
	lookup[561] = -12'sd606;
	lookup[562] = -12'sd618;
	lookup[563] = -12'sd630;
	lookup[564] = -12'sd642;
	lookup[565] = -12'sd654;
	lookup[566] = -12'sd666;
	lookup[567] = -12'sd678;
	lookup[568] = -12'sd689;
	lookup[569] = -12'sd701;
	lookup[570] = -12'sd713;
	lookup[571] = -12'sd725;
	lookup[572] = -12'sd737;
	lookup[573] = -12'sd748;
	lookup[574] = -12'sd760;
	lookup[575] = -12'sd772;
	lookup[576] = -12'sd783;
	lookup[577] = -12'sd795;
	lookup[578] = -12'sd806;
	lookup[579] = -12'sd818;
	lookup[580] = -12'sd829;
	lookup[581] = -12'sd841;
	lookup[582] = -12'sd852;
	lookup[583] = -12'sd864;
	lookup[584] = -12'sd875;
	lookup[585] = -12'sd886;
	lookup[586] = -12'sd898;
	lookup[587] = -12'sd909;
	lookup[588] = -12'sd920;
	lookup[589] = -12'sd932;
	lookup[590] = -12'sd943;
	lookup[591] = -12'sd954;
	lookup[592] = -12'sd965;
	lookup[593] = -12'sd976;
	lookup[594] = -12'sd987;
	lookup[595] = -12'sd998;
	lookup[596] = -12'sd1009;
	lookup[597] = -12'sd1020;
	lookup[598] = -12'sd1031;
	lookup[599] = -12'sd1042;
	lookup[600] = -12'sd1052;
	lookup[601] = -12'sd1063;
	lookup[602] = -12'sd1074;
	lookup[603] = -12'sd1085;
	lookup[604] = -12'sd1095;
	lookup[605] = -12'sd1106;
	lookup[606] = -12'sd1116;
	lookup[607] = -12'sd1127;
	lookup[608] = -12'sd1137;
	lookup[609] = -12'sd1148;
	lookup[610] = -12'sd1158;
	lookup[611] = -12'sd1168;
	lookup[612] = -12'sd1179;
	lookup[613] = -12'sd1189;
	lookup[614] = -12'sd1199;
	lookup[615] = -12'sd1209;
	lookup[616] = -12'sd1219;
	lookup[617] = -12'sd1230;
	lookup[618] = -12'sd1240;
	lookup[619] = -12'sd1250;
	lookup[620] = -12'sd1259;
	lookup[621] = -12'sd1269;
	lookup[622] = -12'sd1279;
	lookup[623] = -12'sd1289;
	lookup[624] = -12'sd1299;
	lookup[625] = -12'sd1308;
	lookup[626] = -12'sd1318;
	lookup[627] = -12'sd1328;
	lookup[628] = -12'sd1337;
	lookup[629] = -12'sd1347;
	lookup[630] = -12'sd1356;
	lookup[631] = -12'sd1366;
	lookup[632] = -12'sd1375;
	lookup[633] = -12'sd1384;
	lookup[634] = -12'sd1393;
	lookup[635] = -12'sd1403;
	lookup[636] = -12'sd1412;
	lookup[637] = -12'sd1421;
	lookup[638] = -12'sd1430;
	lookup[639] = -12'sd1439;
	lookup[640] = -12'sd1448;
	lookup[641] = -12'sd1457;
	lookup[642] = -12'sd1465;
	lookup[643] = -12'sd1474;
	lookup[644] = -12'sd1483;
	lookup[645] = -12'sd1491;
	lookup[646] = -12'sd1500;
	lookup[647] = -12'sd1509;
	lookup[648] = -12'sd1517;
	lookup[649] = -12'sd1525;
	lookup[650] = -12'sd1534;
	lookup[651] = -12'sd1542;
	lookup[652] = -12'sd1550;
	lookup[653] = -12'sd1558;
	lookup[654] = -12'sd1567;
	lookup[655] = -12'sd1575;
	lookup[656] = -12'sd1583;
	lookup[657] = -12'sd1591;
	lookup[658] = -12'sd1598;
	lookup[659] = -12'sd1606;
	lookup[660] = -12'sd1614;
	lookup[661] = -12'sd1622;
	lookup[662] = -12'sd1629;
	lookup[663] = -12'sd1637;
	lookup[664] = -12'sd1644;
	lookup[665] = -12'sd1652;
	lookup[666] = -12'sd1659;
	lookup[667] = -12'sd1667;
	lookup[668] = -12'sd1674;
	lookup[669] = -12'sd1681;
	lookup[670] = -12'sd1688;
	lookup[671] = -12'sd1695;
	lookup[672] = -12'sd1702;
	lookup[673] = -12'sd1709;
	lookup[674] = -12'sd1716;
	lookup[675] = -12'sd1723;
	lookup[676] = -12'sd1730;
	lookup[677] = -12'sd1736;
	lookup[678] = -12'sd1743;
	lookup[679] = -12'sd1750;
	lookup[680] = -12'sd1756;
	lookup[681] = -12'sd1763;
	lookup[682] = -12'sd1769;
	lookup[683] = -12'sd1775;
	lookup[684] = -12'sd1781;
	lookup[685] = -12'sd1788;
	lookup[686] = -12'sd1794;
	lookup[687] = -12'sd1800;
	lookup[688] = -12'sd1806;
	lookup[689] = -12'sd1812;
	lookup[690] = -12'sd1817;
	lookup[691] = -12'sd1823;
	lookup[692] = -12'sd1829;
	lookup[693] = -12'sd1834;
	lookup[694] = -12'sd1840;
	lookup[695] = -12'sd1845;
	lookup[696] = -12'sd1851;
	lookup[697] = -12'sd1856;
	lookup[698] = -12'sd1861;
	lookup[699] = -12'sd1867;
	lookup[700] = -12'sd1872;
	lookup[701] = -12'sd1877;
	lookup[702] = -12'sd1882;
	lookup[703] = -12'sd1887;
	lookup[704] = -12'sd1892;
	lookup[705] = -12'sd1896;
	lookup[706] = -12'sd1901;
	lookup[707] = -12'sd1906;
	lookup[708] = -12'sd1910;
	lookup[709] = -12'sd1915;
	lookup[710] = -12'sd1919;
	lookup[711] = -12'sd1924;
	lookup[712] = -12'sd1928;
	lookup[713] = -12'sd1932;
	lookup[714] = -12'sd1936;
	lookup[715] = -12'sd1940;
	lookup[716] = -12'sd1944;
	lookup[717] = -12'sd1948;
	lookup[718] = -12'sd1952;
	lookup[719] = -12'sd1956;
	lookup[720] = -12'sd1959;
	lookup[721] = -12'sd1963;
	lookup[722] = -12'sd1966;
	lookup[723] = -12'sd1970;
	lookup[724] = -12'sd1973;
	lookup[725] = -12'sd1977;
	lookup[726] = -12'sd1980;
	lookup[727] = -12'sd1983;
	lookup[728] = -12'sd1986;
	lookup[729] = -12'sd1989;
	lookup[730] = -12'sd1992;
	lookup[731] = -12'sd1995;
	lookup[732] = -12'sd1998;
	lookup[733] = -12'sd2000;
	lookup[734] = -12'sd2003;
	lookup[735] = -12'sd2006;
	lookup[736] = -12'sd2008;
	lookup[737] = -12'sd2011;
	lookup[738] = -12'sd2013;
	lookup[739] = -12'sd2015;
	lookup[740] = -12'sd2017;
	lookup[741] = -12'sd2019;
	lookup[742] = -12'sd2021;
	lookup[743] = -12'sd2023;
	lookup[744] = -12'sd2025;
	lookup[745] = -12'sd2027;
	lookup[746] = -12'sd2029;
	lookup[747] = -12'sd2031;
	lookup[748] = -12'sd2032;
	lookup[749] = -12'sd2034;
	lookup[750] = -12'sd2035;
	lookup[751] = -12'sd2036;
	lookup[752] = -12'sd2038;
	lookup[753] = -12'sd2039;
	lookup[754] = -12'sd2040;
	lookup[755] = -12'sd2041;
	lookup[756] = -12'sd2042;
	lookup[757] = -12'sd2043;
	lookup[758] = -12'sd2044;
	lookup[759] = -12'sd2044;
	lookup[760] = -12'sd2045;
	lookup[761] = -12'sd2046;
	lookup[762] = -12'sd2046;
	lookup[763] = -12'sd2047;
	lookup[764] = -12'sd2047;
	lookup[765] = -12'sd2047;
	lookup[766] = -12'sd2047;
	lookup[767] = -12'sd2047;
	lookup[768] = -12'sd2047;
	lookup[769] = -12'sd2047;
	lookup[770] = -12'sd2047;
	lookup[771] = -12'sd2047;
	lookup[772] = -12'sd2047;
	lookup[773] = -12'sd2047;
	lookup[774] = -12'sd2046;
	lookup[775] = -12'sd2046;
	lookup[776] = -12'sd2045;
	lookup[777] = -12'sd2044;
	lookup[778] = -12'sd2044;
	lookup[779] = -12'sd2043;
	lookup[780] = -12'sd2042;
	lookup[781] = -12'sd2041;
	lookup[782] = -12'sd2040;
	lookup[783] = -12'sd2039;
	lookup[784] = -12'sd2038;
	lookup[785] = -12'sd2036;
	lookup[786] = -12'sd2035;
	lookup[787] = -12'sd2034;
	lookup[788] = -12'sd2032;
	lookup[789] = -12'sd2031;
	lookup[790] = -12'sd2029;
	lookup[791] = -12'sd2027;
	lookup[792] = -12'sd2025;
	lookup[793] = -12'sd2023;
	lookup[794] = -12'sd2021;
	lookup[795] = -12'sd2019;
	lookup[796] = -12'sd2017;
	lookup[797] = -12'sd2015;
	lookup[798] = -12'sd2013;
	lookup[799] = -12'sd2011;
	lookup[800] = -12'sd2008;
	lookup[801] = -12'sd2006;
	lookup[802] = -12'sd2003;
	lookup[803] = -12'sd2000;
	lookup[804] = -12'sd1998;
	lookup[805] = -12'sd1995;
	lookup[806] = -12'sd1992;
	lookup[807] = -12'sd1989;
	lookup[808] = -12'sd1986;
	lookup[809] = -12'sd1983;
	lookup[810] = -12'sd1980;
	lookup[811] = -12'sd1977;
	lookup[812] = -12'sd1973;
	lookup[813] = -12'sd1970;
	lookup[814] = -12'sd1966;
	lookup[815] = -12'sd1963;
	lookup[816] = -12'sd1959;
	lookup[817] = -12'sd1956;
	lookup[818] = -12'sd1952;
	lookup[819] = -12'sd1948;
	lookup[820] = -12'sd1944;
	lookup[821] = -12'sd1940;
	lookup[822] = -12'sd1936;
	lookup[823] = -12'sd1932;
	lookup[824] = -12'sd1928;
	lookup[825] = -12'sd1924;
	lookup[826] = -12'sd1919;
	lookup[827] = -12'sd1915;
	lookup[828] = -12'sd1910;
	lookup[829] = -12'sd1906;
	lookup[830] = -12'sd1901;
	lookup[831] = -12'sd1896;
	lookup[832] = -12'sd1892;
	lookup[833] = -12'sd1887;
	lookup[834] = -12'sd1882;
	lookup[835] = -12'sd1877;
	lookup[836] = -12'sd1872;
	lookup[837] = -12'sd1867;
	lookup[838] = -12'sd1861;
	lookup[839] = -12'sd1856;
	lookup[840] = -12'sd1851;
	lookup[841] = -12'sd1845;
	lookup[842] = -12'sd1840;
	lookup[843] = -12'sd1834;
	lookup[844] = -12'sd1829;
	lookup[845] = -12'sd1823;
	lookup[846] = -12'sd1817;
	lookup[847] = -12'sd1812;
	lookup[848] = -12'sd1806;
	lookup[849] = -12'sd1800;
	lookup[850] = -12'sd1794;
	lookup[851] = -12'sd1788;
	lookup[852] = -12'sd1781;
	lookup[853] = -12'sd1775;
	lookup[854] = -12'sd1769;
	lookup[855] = -12'sd1763;
	lookup[856] = -12'sd1756;
	lookup[857] = -12'sd1750;
	lookup[858] = -12'sd1743;
	lookup[859] = -12'sd1736;
	lookup[860] = -12'sd1730;
	lookup[861] = -12'sd1723;
	lookup[862] = -12'sd1716;
	lookup[863] = -12'sd1709;
	lookup[864] = -12'sd1702;
	lookup[865] = -12'sd1695;
	lookup[866] = -12'sd1688;
	lookup[867] = -12'sd1681;
	lookup[868] = -12'sd1674;
	lookup[869] = -12'sd1667;
	lookup[870] = -12'sd1659;
	lookup[871] = -12'sd1652;
	lookup[872] = -12'sd1644;
	lookup[873] = -12'sd1637;
	lookup[874] = -12'sd1629;
	lookup[875] = -12'sd1622;
	lookup[876] = -12'sd1614;
	lookup[877] = -12'sd1606;
	lookup[878] = -12'sd1598;
	lookup[879] = -12'sd1591;
	lookup[880] = -12'sd1583;
	lookup[881] = -12'sd1575;
	lookup[882] = -12'sd1567;
	lookup[883] = -12'sd1558;
	lookup[884] = -12'sd1550;
	lookup[885] = -12'sd1542;
	lookup[886] = -12'sd1534;
	lookup[887] = -12'sd1525;
	lookup[888] = -12'sd1517;
	lookup[889] = -12'sd1509;
	lookup[890] = -12'sd1500;
	lookup[891] = -12'sd1491;
	lookup[892] = -12'sd1483;
	lookup[893] = -12'sd1474;
	lookup[894] = -12'sd1465;
	lookup[895] = -12'sd1457;
	lookup[896] = -12'sd1448;
	lookup[897] = -12'sd1439;
	lookup[898] = -12'sd1430;
	lookup[899] = -12'sd1421;
	lookup[900] = -12'sd1412;
	lookup[901] = -12'sd1403;
	lookup[902] = -12'sd1393;
	lookup[903] = -12'sd1384;
	lookup[904] = -12'sd1375;
	lookup[905] = -12'sd1366;
	lookup[906] = -12'sd1356;
	lookup[907] = -12'sd1347;
	lookup[908] = -12'sd1337;
	lookup[909] = -12'sd1328;
	lookup[910] = -12'sd1318;
	lookup[911] = -12'sd1308;
	lookup[912] = -12'sd1299;
	lookup[913] = -12'sd1289;
	lookup[914] = -12'sd1279;
	lookup[915] = -12'sd1269;
	lookup[916] = -12'sd1259;
	lookup[917] = -12'sd1250;
	lookup[918] = -12'sd1240;
	lookup[919] = -12'sd1230;
	lookup[920] = -12'sd1219;
	lookup[921] = -12'sd1209;
	lookup[922] = -12'sd1199;
	lookup[923] = -12'sd1189;
	lookup[924] = -12'sd1179;
	lookup[925] = -12'sd1168;
	lookup[926] = -12'sd1158;
	lookup[927] = -12'sd1148;
	lookup[928] = -12'sd1137;
	lookup[929] = -12'sd1127;
	lookup[930] = -12'sd1116;
	lookup[931] = -12'sd1106;
	lookup[932] = -12'sd1095;
	lookup[933] = -12'sd1085;
	lookup[934] = -12'sd1074;
	lookup[935] = -12'sd1063;
	lookup[936] = -12'sd1052;
	lookup[937] = -12'sd1042;
	lookup[938] = -12'sd1031;
	lookup[939] = -12'sd1020;
	lookup[940] = -12'sd1009;
	lookup[941] = -12'sd998;
	lookup[942] = -12'sd987;
	lookup[943] = -12'sd976;
	lookup[944] = -12'sd965;
	lookup[945] = -12'sd954;
	lookup[946] = -12'sd943;
	lookup[947] = -12'sd932;
	lookup[948] = -12'sd920;
	lookup[949] = -12'sd909;
	lookup[950] = -12'sd898;
	lookup[951] = -12'sd886;
	lookup[952] = -12'sd875;
	lookup[953] = -12'sd864;
	lookup[954] = -12'sd852;
	lookup[955] = -12'sd841;
	lookup[956] = -12'sd829;
	lookup[957] = -12'sd818;
	lookup[958] = -12'sd806;
	lookup[959] = -12'sd795;
	lookup[960] = -12'sd783;
	lookup[961] = -12'sd772;
	lookup[962] = -12'sd760;
	lookup[963] = -12'sd748;
	lookup[964] = -12'sd737;
	lookup[965] = -12'sd725;
	lookup[966] = -12'sd713;
	lookup[967] = -12'sd701;
	lookup[968] = -12'sd689;
	lookup[969] = -12'sd678;
	lookup[970] = -12'sd666;
	lookup[971] = -12'sd654;
	lookup[972] = -12'sd642;
	lookup[973] = -12'sd630;
	lookup[974] = -12'sd618;
	lookup[975] = -12'sd606;
	lookup[976] = -12'sd594;
	lookup[977] = -12'sd582;
	lookup[978] = -12'sd570;
	lookup[979] = -12'sd558;
	lookup[980] = -12'sd546;
	lookup[981] = -12'sd534;
	lookup[982] = -12'sd521;
	lookup[983] = -12'sd509;
	lookup[984] = -12'sd497;
	lookup[985] = -12'sd485;
	lookup[986] = -12'sd473;
	lookup[987] = -12'sd460;
	lookup[988] = -12'sd448;
	lookup[989] = -12'sd436;
	lookup[990] = -12'sd424;
	lookup[991] = -12'sd411;
	lookup[992] = -12'sd399;
	lookup[993] = -12'sd387;
	lookup[994] = -12'sd374;
	lookup[995] = -12'sd362;
	lookup[996] = -12'sd350;
	lookup[997] = -12'sd337;
	lookup[998] = -12'sd325;
	lookup[999] = -12'sd312;
	lookup[1000] = -12'sd300;
	lookup[1001] = -12'sd288;
	lookup[1002] = -12'sd275;
	lookup[1003] = -12'sd263;
	lookup[1004] = -12'sd250;
	lookup[1005] = -12'sd238;
	lookup[1006] = -12'sd225;
	lookup[1007] = -12'sd213;
	lookup[1008] = -12'sd200;
	lookup[1009] = -12'sd188;
	lookup[1010] = -12'sd175;
	lookup[1011] = -12'sd163;
	lookup[1012] = -12'sd150;
	lookup[1013] = -12'sd138;
	lookup[1014] = -12'sd125;
	lookup[1015] = -12'sd113;
	lookup[1016] = -12'sd100;
	lookup[1017] = -12'sd87;
	lookup[1018] = -12'sd75;
	lookup[1019] = -12'sd62;
	lookup[1020] = -12'sd50;
	lookup[1021] = -12'sd37;
	lookup[1022] = -12'sd25;
	lookup[1023] = -12'sd12;
end


endmodule
